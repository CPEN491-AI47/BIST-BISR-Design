`define WORD_SIZE 16
`define ROWS 2
`define COLS 2 
`define ENABLE_RANDOM
`define SEED 100
`define ENABLE_FI
`define ENABLE_TMR