`define WORD_SIZE 16
`define ROWS 2
`define COLS 2 
`define SEED 100

`define stw_mult_op1 4
`define stw_mult_op2 3
`define stw_add_op 1
`define stw_expected_out 13
// `define ENABLE_RANDOM
// `define ENABLE_TMR

`define ENABLE_FI
`define ENABLE_STW
`define ENABLE_WPROXY