`define WORD_SIZE 16
`define ROWS 3
`define COLS 3 
`define SEED 100
// `define ENABLE_RANDOM
// `define ENABLE_TMR

`define ENABLE_FI
`define ENABLE_STW
`define ENABLE_WPROXY